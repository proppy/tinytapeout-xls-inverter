module user_module_USER_MODULE_ID(
  input wire [7:0] io_in,
  output wire [7:0] out
);
  assign out = ~io_in;
endmodule
